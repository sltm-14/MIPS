/******************************************************************
* Description
*		This is an AND gate:
*
******************************************************************/
module ANDGate
(
	input A,
	input B,

	output C
);


	assign C = A & B;

endmodule
