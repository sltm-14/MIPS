/******************************************************************
* Description
*	This a file to include all the definitions needed in the compilation process
*
******************************************************************/

/*If this constant is defined, it allows to include sentences that are used in the simulation
*  process in modelsim. If it is not defined, it allows to synthesize the processor in Quartus II.
* In order to undefine the constant, it must be commented. Note that the apostrophe is part of the definition*/

//`define MONITORS //Constant definitions

module Definitions(

    );

endmodule
