/******************************************************************
* Description
*		OR gate
*
******************************************************************/
module OR_Gate
(
	input  A,
	input  B,

	output C
);

	assign C = A | B;

endmodule
