library verilog;
use verilog.vl_types.all;
entity Definitions is
end Definitions;
